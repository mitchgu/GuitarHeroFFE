module SC_buffer_serializer(
    input clk,
    input song_time,
    input [36:0] match_trigger,
    input [37*16-1:0] match_time
    
    
    
    );
    
    
endmodule