module AV_block(
    
    
    
    
    );
    
endmodule