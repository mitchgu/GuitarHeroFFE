module AV_note_sprite(
    input clk65,
    input [10:0] x,
    input [9:0] y,
    input [10:0] hcount,
    input [9:0] vcount,
    input [4:0] value,
    
    output reg [12:0] note_pixel
    
    );
    
    
    
    
    
    initial note_pixel <= 0;
    
    
    
endmodule