module SC_score(
    input clk, //100mhz clk
    input [15:0] dt, //margin of correctness for a matched note
    input en, //match enable
    
    output reg score //total score DETERMINE WIDTH
    );
    
    
    
    
    
    
    
endmodule