module SC_note_matching_super(
    input clk,
    input [36:0] NDATA,
    
    
    
    );
    
    reg [36:0] note_prev; //array of previous note-states
    
    
    
    
endmodule