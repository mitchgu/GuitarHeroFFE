module CL_block(
    
    
    
    
    
    );
    
    
endmodule