`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:54:30 10/28/2014 
// Design Name: 
// Module Name:    pwm_module 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module pwm11 ( 
    input clk,
    input [10:0] PWM_in, 
    output reg PWM_out,
    output PWM_sd
    );

    reg [10:0] new_pwm=0;
    reg [10:0] PWM_ramp=0; 
    always @(posedge clk) begin
        if (PWM_ramp==0) new_pwm <= PWM_in;
        PWM_ramp <= PWM_ramp + 1'b1;
        PWM_out <= (new_pwm>PWM_ramp);
    end

    assign PWM_sd = 1;

endmodule