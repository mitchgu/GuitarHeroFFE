module SC_block(
    
    
    
    
    
    
    
    );
    
    
    
endmodule